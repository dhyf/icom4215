module main;
  initial 
    begin
      $display("Hello");
      $finish ;
    end
endmodule
